

module sine_gen(
	input	wire	clk,
	input 	wire 	rst,
	input   wire	send,
	output  wire	[15:0]  sine
    );

reg [15:0]  q;
reg [9:0]   ms; // main state

assign sine = q;

localparam
    ms_pause    = 10'd0,
    ms_1        = 10'd1,
    ms_2        = 10'd2,
    ms_3        = 10'd3,
    ms_4        = 10'd4,
    ms_5        = 10'd5,
    ms_6        = 10'd6,
    ms_7        = 10'd7,
    ms_8        = 10'd8,
    ms_9        = 10'd9,
    ms_10        = 10'd10,
    ms_11        = 10'd11,
    ms_12        = 10'd12,
    ms_13        = 10'd13,
    ms_14        = 10'd14,
    ms_15        = 10'd15,
    ms_16        = 10'd16,
    ms_17        = 10'd17,
    ms_18        = 10'd18,
    ms_19        = 10'd19,
    ms_20        = 10'd20,
    ms_21        = 10'd21,
    ms_22        = 10'd22,
    ms_23        = 10'd23,
    ms_24        = 10'd24,
    ms_25        = 10'd25,
    ms_26        = 10'd26,
    ms_27        = 10'd27,
    ms_28        = 10'd28,
    ms_29        = 10'd29,
    ms_30        = 10'd30,
    ms_31        = 10'd31,
    ms_32        = 10'd32,
    ms_33        = 10'd33,
    ms_34        = 10'd34,
    ms_35        = 10'd35,
    ms_36        = 10'd36,
    ms_37        = 10'd37,
    ms_38        = 10'd38,
    ms_39        = 10'd39,
    ms_40        = 10'd40,
    ms_41        = 10'd41,
    ms_42        = 10'd42,
    ms_43        = 10'd43,
    ms_44        = 10'd44,
    ms_45        = 10'd45,
    ms_46        = 10'd46,
    ms_47        = 10'd47,
    ms_48        = 10'd48,
    ms_49        = 10'd49,
    ms_50        = 10'd50,
    ms_51        = 10'd51,
    ms_52        = 10'd52,
    ms_53        = 10'd53,
    ms_54        = 10'd54,
    ms_55        = 10'd55,
    ms_56        = 10'd56,
    ms_57        = 10'd57,
    ms_58        = 10'd58,
    ms_59        = 10'd59,
    ms_60        = 10'd60,
    ms_61        = 10'd61,
    ms_62        = 10'd62,
    ms_63        = 10'd63,
    ms_64        = 10'd64,
    ms_65        = 10'd65,
    ms_66        = 10'd66,
    ms_67        = 10'd67,
    ms_68        = 10'd68,
    ms_69        = 10'd69,
    ms_70        = 10'd70,
    ms_71        = 10'd71,
    ms_72        = 10'd72,
    ms_73        = 10'd73,
    ms_74        = 10'd74,
    ms_75        = 10'd75,
    ms_76        = 10'd76,
    ms_77        = 10'd77,
    ms_78        = 10'd78,
    ms_79        = 10'd79,
    ms_80        = 10'd80,
    ms_81        = 10'd81,
    ms_82        = 10'd82,
    ms_83        = 10'd83,
    ms_84        = 10'd84,
    ms_85        = 10'd85,
    ms_86        = 10'd86,
    ms_87        = 10'd87,
    ms_88        = 10'd88,
    ms_89        = 10'd89,
    ms_90        = 10'd90,
    ms_91        = 10'd91,
    ms_92        = 10'd92,
    ms_93        = 10'd93,
    ms_94        = 10'd94,
    ms_95        = 10'd95,
    ms_96        = 10'd96,
    ms_97        = 10'd97,
    ms_98        = 10'd98,
    ms_99        = 10'd99,
    ms_100        = 10'd100,
    ms_101        = 10'd101,
    ms_102        = 10'd102,
    ms_103        = 10'd103,
    ms_104        = 10'd104,
    ms_105        = 10'd105,
    ms_106        = 10'd106,
    ms_107        = 10'd107,
    ms_108        = 10'd108,
    ms_109        = 10'd109,
    ms_110        = 10'd110,
    ms_111        = 10'd111,
    ms_112        = 10'd112,
    ms_113        = 10'd113,
    ms_114        = 10'd114,
    ms_115        = 10'd115,
    ms_116        = 10'd116,
    ms_117        = 10'd117,
    ms_118        = 10'd118,
    ms_119        = 10'd119,
    ms_120        = 10'd120,
    ms_121        = 10'd121,
    ms_122        = 10'd122,
    ms_123        = 10'd123,
    ms_124        = 10'd124,
    ms_125        = 10'd125,
    ms_126        = 10'd126,
    ms_127        = 10'd127,
    ms_128        = 10'd128,
    ms_129        = 10'd129,
    ms_130        = 10'd130,
    ms_131        = 10'd131,
    ms_132        = 10'd132,
    ms_133        = 10'd133,
    ms_134        = 10'd134,
    ms_135        = 10'd135,
    ms_136        = 10'd136,
    ms_137        = 10'd137,
    ms_138        = 10'd138,
    ms_139        = 10'd139,
    ms_140        = 10'd140,
    ms_141        = 10'd141,
    ms_142        = 10'd142,
    ms_143        = 10'd143,
    ms_144        = 10'd144,
    ms_145        = 10'd145,
    ms_146        = 10'd146,
    ms_147        = 10'd147,
    ms_148        = 10'd148,
    ms_149        = 10'd149,
    ms_150        = 10'd150,
    ms_151        = 10'd151,
    ms_152        = 10'd152,
    ms_153        = 10'd153,
    ms_154        = 10'd154,
    ms_155        = 10'd155,
    ms_156        = 10'd156,
    ms_157        = 10'd157,
    ms_158        = 10'd158,
    ms_159        = 10'd159,
    ms_160        = 10'd160,
    ms_161        = 10'd161,
    ms_162        = 10'd162,
    ms_163        = 10'd163,
    ms_164        = 10'd164,
    ms_165        = 10'd165,
    ms_166        = 10'd166,
    ms_167        = 10'd167,
    ms_168        = 10'd168,
    ms_169        = 10'd169,
    ms_170        = 10'd170,
    ms_171        = 10'd171,
    ms_172        = 10'd172,
    ms_173        = 10'd173,
    ms_174        = 10'd174,
    ms_175        = 10'd175,
    ms_176        = 10'd176,
    ms_177        = 10'd177,
    ms_178        = 10'd178,
    ms_179        = 10'd179,
    ms_180        = 10'd180,
    ms_181        = 10'd181,
    ms_182        = 10'd182,
    ms_183        = 10'd183,
    ms_184        = 10'd184,
    ms_185        = 10'd185,
    ms_186        = 10'd186,
    ms_187        = 10'd187,
    ms_188        = 10'd188,
    ms_189        = 10'd189,
    ms_190        = 10'd190,
    ms_191        = 10'd191,
    ms_192        = 10'd192,
    ms_193        = 10'd193,
    ms_194        = 10'd194,
    ms_195        = 10'd195,
    ms_196        = 10'd196,
    ms_197        = 10'd197,
    ms_198        = 10'd198,
    ms_199        = 10'd199,
    ms_200        = 10'd200,
    ms_201        = 10'd201,
    ms_202        = 10'd202,
    ms_203        = 10'd203,
    ms_204        = 10'd204,
    ms_205        = 10'd205,
    ms_206        = 10'd206,
    ms_207        = 10'd207,
    ms_208        = 10'd208,
    ms_209        = 10'd209,
    ms_210        = 10'd210,
    ms_211        = 10'd211,
    ms_212        = 10'd212,
    ms_213        = 10'd213,
    ms_214        = 10'd214,
    ms_215        = 10'd215,
    ms_216        = 10'd216,
    ms_217        = 10'd217,
    ms_218        = 10'd218,
    ms_219        = 10'd219,
    ms_220        = 10'd220,
    ms_221        = 10'd221,
    ms_222        = 10'd222,
    ms_223        = 10'd223,
    ms_224        = 10'd224,
    ms_225        = 10'd225,
    ms_226        = 10'd226,
    ms_227        = 10'd227,
    ms_228        = 10'd228,
    ms_229        = 10'd229,
    ms_230        = 10'd230,
    ms_231        = 10'd231,
    ms_232        = 10'd232,
    ms_233        = 10'd233,
    ms_234        = 10'd234,
    ms_235        = 10'd235,
    ms_236        = 10'd236,
    ms_237        = 10'd237,
    ms_238        = 10'd238,
    ms_239        = 10'd239,
    ms_240        = 10'd240,
    ms_241        = 10'd241,
    ms_242        = 10'd242,
    ms_243        = 10'd243,
    ms_244        = 10'd244,
    ms_245        = 10'd245,
    ms_246        = 10'd246,
    ms_247        = 10'd247,
    ms_248        = 10'd248,
    ms_249        = 10'd249,
    ms_250        = 10'd250,
    ms_251        = 10'd251,
    ms_252        = 10'd252,
    ms_253        = 10'd253,
    ms_254        = 10'd254,
    ms_255        = 10'd255,
    ms_256        = 10'd256,
    ms_257        = 10'd257,
    ms_258        = 10'd258,
    ms_259        = 10'd259,
    ms_260        = 10'd260,
    ms_261        = 10'd261,
    ms_262        = 10'd262,
    ms_263        = 10'd263,
    ms_264        = 10'd264,
    ms_265        = 10'd265,
    ms_266        = 10'd266,
    ms_267        = 10'd267,
    ms_268        = 10'd268,
    ms_269        = 10'd269,
    ms_270        = 10'd270,
    ms_271        = 10'd271,
    ms_272        = 10'd272,
    ms_273        = 10'd273,
    ms_274        = 10'd274,
    ms_275        = 10'd275,
    ms_276        = 10'd276,
    ms_277        = 10'd277,
    ms_278        = 10'd278,
    ms_279        = 10'd279,
    ms_280        = 10'd280,
    ms_281        = 10'd281,
    ms_282        = 10'd282,
    ms_283        = 10'd283,
    ms_284        = 10'd284,
    ms_285        = 10'd285,
    ms_286        = 10'd286,
    ms_287        = 10'd287,
    ms_288        = 10'd288,
    ms_289        = 10'd289,
    ms_290        = 10'd290,
    ms_291        = 10'd291,
    ms_292        = 10'd292,
    ms_293        = 10'd293,
    ms_294        = 10'd294,
    ms_295        = 10'd295,
    ms_296        = 10'd296,
    ms_297        = 10'd297,
    ms_298        = 10'd298,
    ms_299        = 10'd299,
    ms_300        = 10'd300,
    ms_301        = 10'd301,
    ms_302        = 10'd302,
    ms_303        = 10'd303,
    ms_304        = 10'd304,
    ms_305        = 10'd305,
    ms_306        = 10'd306,
    ms_307        = 10'd307,
    ms_308        = 10'd308,
    ms_309        = 10'd309,
    ms_310        = 10'd310,
    ms_311        = 10'd311,
    ms_312        = 10'd312,
    ms_313        = 10'd313,
    ms_314        = 10'd314,
    ms_315        = 10'd315,
    ms_316        = 10'd316,
    ms_317        = 10'd317,
    ms_318        = 10'd318,
    ms_319        = 10'd319,
    ms_320        = 10'd320,
    ms_321        = 10'd321,
    ms_322        = 10'd322,
    ms_323        = 10'd323,
    ms_324        = 10'd324,
    ms_325        = 10'd325,
    ms_326        = 10'd326,
    ms_327        = 10'd327,
    ms_328        = 10'd328,
    ms_329        = 10'd329,
    ms_330        = 10'd330,
    ms_331        = 10'd331,
    ms_332        = 10'd332,
    ms_333        = 10'd333,
    ms_334        = 10'd334,
    ms_335        = 10'd335,
    ms_336        = 10'd336,
    ms_337        = 10'd337,
    ms_338        = 10'd338,
    ms_339        = 10'd339,
    ms_340        = 10'd340,
    ms_341        = 10'd341,
    ms_342        = 10'd342,
    ms_343        = 10'd343,
    ms_344        = 10'd344,
    ms_345        = 10'd345,
    ms_346        = 10'd346,
    ms_347        = 10'd347,
    ms_348        = 10'd348,
    ms_349        = 10'd349,
    ms_350        = 10'd350,
    ms_351        = 10'd351,
    ms_352        = 10'd352,
    ms_353        = 10'd353,
    ms_354        = 10'd354,
    ms_355        = 10'd355,
    ms_356        = 10'd356,
    ms_357        = 10'd357,
    ms_358        = 10'd358,
    ms_359        = 10'd359,
    ms_360        = 10'd360,
    ms_361        = 10'd361,
    ms_362        = 10'd362,
    ms_363        = 10'd363,
    ms_364        = 10'd364,
    ms_365        = 10'd365,
    ms_366        = 10'd366,
    ms_367        = 10'd367,
    ms_368        = 10'd368,
    ms_369        = 10'd369,
    ms_370        = 10'd370,
    ms_371        = 10'd371,
    ms_372        = 10'd372,
    ms_373        = 10'd373,
    ms_374        = 10'd374,
    ms_375        = 10'd375,
    ms_376        = 10'd376,
    ms_377        = 10'd377,
    ms_378        = 10'd378,
    ms_379        = 10'd379,
    ms_380        = 10'd380,
    ms_381        = 10'd381,
    ms_382        = 10'd382,
    ms_383        = 10'd383,
    ms_384        = 10'd384,
    ms_385        = 10'd385,
    ms_386        = 10'd386,
    ms_387        = 10'd387,
    ms_388        = 10'd388,
    ms_389        = 10'd389,
    ms_390        = 10'd390,
    ms_391        = 10'd391,
    ms_392        = 10'd392,
    ms_393        = 10'd393,
    ms_394        = 10'd394,
    ms_395        = 10'd395,
    ms_396        = 10'd396,
    ms_397        = 10'd397,
    ms_398        = 10'd398,
    ms_399        = 10'd399,
    ms_400        = 10'd400,
    ms_401        = 10'd401,
    ms_402        = 10'd402,
    ms_403        = 10'd403,
    ms_404        = 10'd404,
    ms_405        = 10'd405,
    ms_406        = 10'd406,
    ms_407        = 10'd407,
    ms_408        = 10'd408,
    ms_409        = 10'd409,
    ms_410        = 10'd410,
    ms_411        = 10'd411,
    ms_412        = 10'd412,
    ms_413        = 10'd413,
    ms_414        = 10'd414,
    ms_415        = 10'd415,
    ms_416        = 10'd416,
    ms_417        = 10'd417,
    ms_418        = 10'd418,
    ms_419        = 10'd419,
    ms_420        = 10'd420,
    ms_421        = 10'd421,
    ms_422        = 10'd422,
    ms_423        = 10'd423,
    ms_424        = 10'd424,
    ms_425        = 10'd425,
    ms_426        = 10'd426,
    ms_427        = 10'd427,
    ms_428        = 10'd428,
    ms_429        = 10'd429,
    ms_430        = 10'd430,
    ms_431        = 10'd431,
    ms_432        = 10'd432,
    ms_433        = 10'd433,
    ms_434        = 10'd434,
    ms_435        = 10'd435,
    ms_436        = 10'd436,
    ms_437        = 10'd437,
    ms_438        = 10'd438,
    ms_439        = 10'd439,
    ms_440        = 10'd440,
    ms_441        = 10'd441,
    ms_442        = 10'd442,
    ms_443        = 10'd443,
    ms_444        = 10'd444,
    ms_445        = 10'd445,
    ms_446        = 10'd446,
    ms_447        = 10'd447,
    ms_448        = 10'd448,
    ms_449        = 10'd449,
    ms_450        = 10'd450,
    ms_451        = 10'd451,
    ms_452        = 10'd452,
    ms_453        = 10'd453,
    ms_454        = 10'd454,
    ms_455        = 10'd455,
    ms_456        = 10'd456,
    ms_457        = 10'd457,
    ms_458        = 10'd458,
    ms_459        = 10'd459,
    ms_460        = 10'd460,
    ms_461        = 10'd461,
    ms_462        = 10'd462,
    ms_463        = 10'd463,
    ms_464        = 10'd464,
    ms_465        = 10'd465,
    ms_466        = 10'd466,
    ms_467        = 10'd467,
    ms_468        = 10'd468,
    ms_469        = 10'd469,
    ms_470        = 10'd470,
    ms_471        = 10'd471,
    ms_472        = 10'd472,
    ms_473        = 10'd473,
    ms_474        = 10'd474,
    ms_475        = 10'd475,
    ms_476        = 10'd476,
    ms_477        = 10'd477,
    ms_478        = 10'd478,
    ms_479        = 10'd479,
    ms_480        = 10'd480,
    ms_481        = 10'd481,
    ms_482        = 10'd482,
    ms_483        = 10'd483,
    ms_484        = 10'd484,
    ms_485        = 10'd485,
    ms_486        = 10'd486,
    ms_487        = 10'd487,
    ms_488        = 10'd488,
    ms_489        = 10'd489,
    ms_490        = 10'd490,
    ms_491        = 10'd491,
    ms_492        = 10'd492,
    ms_493        = 10'd493,
    ms_494        = 10'd494,
    ms_495        = 10'd495,
    ms_496        = 10'd496,
    ms_497        = 10'd497,
    ms_498        = 10'd498,
    ms_499        = 10'd499,
    ms_500        = 10'd500,
    ms_501        = 10'd501,
    ms_502        = 10'd502,
    ms_503        = 10'd503,
    ms_504        = 10'd504,
    ms_505        = 10'd505,
    ms_506        = 10'd506,
    ms_507        = 10'd507,
    ms_508        = 10'd508,
    ms_509        = 10'd509,
    ms_510        = 10'd510,
    ms_511        = 10'd511,
    ms_512        = 10'd512,
    ms_513        = 10'd513,
    ms_514        = 10'd514,
    ms_515        = 10'd515,
    ms_516        = 10'd516,
    ms_517        = 10'd517,
    ms_518        = 10'd518,
    ms_519        = 10'd519,
    ms_520        = 10'd520,
    ms_521        = 10'd521,
    ms_522        = 10'd522,
    ms_523        = 10'd523,
    ms_524        = 10'd524,
    ms_525        = 10'd525,
    ms_526        = 10'd526,
    ms_527        = 10'd527,
    ms_528        = 10'd528,
    ms_529        = 10'd529,
    ms_530        = 10'd530,
    ms_531        = 10'd531,
    ms_532        = 10'd532,
    ms_533        = 10'd533,
    ms_534        = 10'd534,
    ms_535        = 10'd535,
    ms_536        = 10'd536,
    ms_537        = 10'd537,
    ms_538        = 10'd538,
    ms_539        = 10'd539,
    ms_540        = 10'd540,
    ms_541        = 10'd541,
    ms_542        = 10'd542,
    ms_543        = 10'd543,
    ms_544        = 10'd544,
    ms_545        = 10'd545,
    ms_546        = 10'd546,
    ms_547        = 10'd547,
    ms_548        = 10'd548,
    ms_549        = 10'd549,
    ms_550        = 10'd550,
    ms_551        = 10'd551,
    ms_552        = 10'd552,
    ms_553        = 10'd553,
    ms_554        = 10'd554,
    ms_555        = 10'd555,
    ms_556        = 10'd556,
    ms_557        = 10'd557,
    ms_558        = 10'd558,
    ms_559        = 10'd559,
    ms_560        = 10'd560,
    ms_561        = 10'd561,
    ms_562        = 10'd562,
    ms_563        = 10'd563,
    ms_564        = 10'd564,
    ms_565        = 10'd565,
    ms_566        = 10'd566,
    ms_567        = 10'd567,
    ms_568        = 10'd568,
    ms_569        = 10'd569,
    ms_570        = 10'd570,
    ms_571        = 10'd571,
    ms_572        = 10'd572,
    ms_573        = 10'd573,
    ms_574        = 10'd574,
    ms_575        = 10'd575,
    ms_576        = 10'd576,
    ms_577        = 10'd577,
    ms_578        = 10'd578,
    ms_579        = 10'd579,
    ms_580        = 10'd580,
    ms_581        = 10'd581,
    ms_582        = 10'd582,
    ms_583        = 10'd583,
    ms_584        = 10'd584,
    ms_585        = 10'd585,
    ms_586        = 10'd586,
    ms_587        = 10'd587,
    ms_588        = 10'd588,
    ms_589        = 10'd589,
    ms_590        = 10'd590,
    ms_591        = 10'd591,
    ms_592        = 10'd592,
    ms_593        = 10'd593,
    ms_594        = 10'd594,
    ms_595        = 10'd595,
    ms_596        = 10'd596,
    ms_597        = 10'd597,
    ms_598        = 10'd598,
    ms_599        = 10'd599,
    ms_600        = 10'd600,
    ms_601        = 10'd601,
    ms_602        = 10'd602,
    ms_603        = 10'd603,
    ms_604        = 10'd604,
    ms_605        = 10'd605,
    ms_606        = 10'd606,
    ms_607        = 10'd607,
    ms_608        = 10'd608,
    ms_609        = 10'd609,
    ms_610        = 10'd610,
    ms_611        = 10'd611,
    ms_612        = 10'd612,
    ms_613        = 10'd613,
    ms_614        = 10'd614,
    ms_615        = 10'd615,
    ms_616        = 10'd616,
    ms_617        = 10'd617,
    ms_618        = 10'd618,
    ms_619        = 10'd619,
    ms_620        = 10'd620,
    ms_621        = 10'd621,
    ms_622        = 10'd622,
    ms_623        = 10'd623,
    ms_624        = 10'd624,
    ms_625        = 10'd625,
    ms_626        = 10'd626,
    ms_627        = 10'd627,
    ms_628        = 10'd628,
    ms_629        = 10'd629,
    ms_630        = 10'd630,
    ms_631        = 10'd631,
    ms_632        = 10'd632,
    ms_633        = 10'd633,
    ms_634        = 10'd634,
    ms_635        = 10'd635,
    ms_636        = 10'd636,
    ms_637        = 10'd637,
    ms_638        = 10'd638,
    ms_639        = 10'd639,
    ms_640        = 10'd640,
    ms_641        = 10'd641,
    ms_642        = 10'd642,
    ms_643        = 10'd643,
    ms_644        = 10'd644,
    ms_645        = 10'd645,
    ms_646        = 10'd646,
    ms_647        = 10'd647,
    ms_648        = 10'd648,
    ms_649        = 10'd649,
    ms_650        = 10'd650,
    ms_651        = 10'd651,
    ms_652        = 10'd652,
    ms_653        = 10'd653,
    ms_654        = 10'd654,
    ms_655        = 10'd655,
    ms_656        = 10'd656,
    ms_657        = 10'd657,
    ms_658        = 10'd658,
    ms_659        = 10'd659,
    ms_660        = 10'd660,
    ms_661        = 10'd661,
    ms_662        = 10'd662,
    ms_663        = 10'd663,
    ms_664        = 10'd664,
    ms_665        = 10'd665,
    ms_666        = 10'd666,
    ms_667        = 10'd667,
    ms_668        = 10'd668,
    ms_669        = 10'd669,
    ms_670        = 10'd670,
    ms_671        = 10'd671,
    ms_672        = 10'd672,
    ms_673        = 10'd673,
    ms_674        = 10'd674,
    ms_675        = 10'd675,
    ms_676        = 10'd676,
    ms_677        = 10'd677,
    ms_678        = 10'd678,
    ms_679        = 10'd679,
    ms_680        = 10'd680,
    ms_681        = 10'd681,
    ms_682        = 10'd682,
    ms_683        = 10'd683,
    ms_684        = 10'd684,
    ms_685        = 10'd685,
    ms_686        = 10'd686,
    ms_687        = 10'd687,
    ms_688        = 10'd688,
    ms_689        = 10'd689,
    ms_690        = 10'd690,
    ms_691        = 10'd691,
    ms_692        = 10'd692,
    ms_693        = 10'd693,
    ms_694        = 10'd694,
    ms_695        = 10'd695,
    ms_696        = 10'd696,
    ms_697        = 10'd697,
    ms_698        = 10'd698,
    ms_699        = 10'd699,
    ms_700        = 10'd700,
    ms_701        = 10'd701,
    ms_702        = 10'd702,
    ms_703        = 10'd703,
    ms_704        = 10'd704,
    ms_705        = 10'd705,
    ms_706        = 10'd706,
    ms_707        = 10'd707,
    ms_708        = 10'd708,
    ms_709        = 10'd709,
    ms_710        = 10'd710,
    ms_711        = 10'd711,
    ms_712        = 10'd712,
    ms_713        = 10'd713,
    ms_714        = 10'd714,
    ms_715        = 10'd715,
    ms_716        = 10'd716,
    ms_717        = 10'd717,
    ms_718        = 10'd718,
    ms_719        = 10'd719,
    ms_720        = 10'd720,
    ms_721        = 10'd721,
    ms_722        = 10'd722,
    ms_723        = 10'd723,
    ms_724        = 10'd724,
    ms_725        = 10'd725,
    ms_726        = 10'd726,
    ms_727        = 10'd727,
    ms_728        = 10'd728,
    ms_729        = 10'd729,
    ms_730        = 10'd730,
    ms_731        = 10'd731,
    ms_732        = 10'd732,
    ms_733        = 10'd733,
    ms_734        = 10'd734,
    ms_735        = 10'd735,
    ms_736        = 10'd736,
    ms_737        = 10'd737,
    ms_738        = 10'd738,
    ms_739        = 10'd739,
    ms_740        = 10'd740,
    ms_741        = 10'd741,
    ms_742        = 10'd742,
    ms_743        = 10'd743,
    ms_744        = 10'd744,
    ms_745        = 10'd745,
    ms_746        = 10'd746,
    ms_747        = 10'd747,
    ms_748        = 10'd748,
    ms_749        = 10'd749,
    ms_750        = 10'd750,
    ms_751        = 10'd751,
    ms_752        = 10'd752,
    ms_753        = 10'd753,
    ms_754        = 10'd754,
    ms_755        = 10'd755,
    ms_756        = 10'd756,
    ms_757        = 10'd757,
    ms_758        = 10'd758,
    ms_759        = 10'd759,
    ms_760        = 10'd760,
    ms_761        = 10'd761,
    ms_762        = 10'd762,
    ms_763        = 10'd763,
    ms_764        = 10'd764,
    ms_765        = 10'd765,
    ms_766        = 10'd766,
    ms_767        = 10'd767,
    ms_768        = 10'd768,
    ms_769        = 10'd769,
    ms_770        = 10'd770,
    ms_771        = 10'd771,
    ms_772        = 10'd772,
    ms_773        = 10'd773,
    ms_774        = 10'd774,
    ms_775        = 10'd775,
    ms_776        = 10'd776,
    ms_777        = 10'd777,
    ms_778        = 10'd778,
    ms_779        = 10'd779,
    ms_780        = 10'd780,
    ms_781        = 10'd781,
    ms_782        = 10'd782,
    ms_783        = 10'd783,
    ms_784        = 10'd784,
    ms_785        = 10'd785,
    ms_786        = 10'd786,
    ms_787        = 10'd787,
    ms_788        = 10'd788,
    ms_789        = 10'd789,
    ms_790        = 10'd790,
    ms_791        = 10'd791,
    ms_792        = 10'd792,
    ms_793        = 10'd793,
    ms_794        = 10'd794,
    ms_795        = 10'd795,
    ms_796        = 10'd796,
    ms_797        = 10'd797,
    ms_798        = 10'd798,
    ms_799        = 10'd799,
    ms_800        = 10'd800;

initial begin
	q <= 16'h8000;
	ms <= ms_pause;
end

always @(posedge rst or posedge clk) begin
	if (rst) begin
		q <= 16'h8000;
		ms <= ms_pause;
	end else begin
	    case (ms) 
		ms_pause: begin
		    q <= 16'h8000;
		    if (send) begin
		        ms <= ms_1;
		    end else begin
		        ms <= ms_pause;
		    end
		end
		ms_1: begin
		    q <= 16'h8000;
		    ms <= ms_2;
		end
		ms_2: begin
		    q <= 16'h8005;
		    ms <= ms_3;
		end
		ms_3: begin
		    q <= 16'h800a;
		    ms <= ms_4;
		end
		ms_4: begin
		    q <= 16'h800f;
		    ms <= ms_5;
		end
		ms_5: begin
		    q <= 16'h8015;
		    ms <= ms_6;
		end
		ms_6: begin
		    q <= 16'h801a;
		    ms <= ms_7;
		end
		ms_7: begin
		    q <= 16'h801f;
		    ms <= ms_8;
		end
		ms_8: begin
		    q <= 16'h8024;
		    ms <= ms_9;
		end
		ms_9: begin
		    q <= 16'h8029;
		    ms <= ms_10;
		end
		ms_10: begin
		    q <= 16'h802e;
		    ms <= ms_11;
		end
		ms_11: begin
		    q <= 16'h8033;
		    ms <= ms_12;
		end
		ms_12: begin
		    q <= 16'h8039;
		    ms <= ms_13;
		end
		ms_13: begin
		    q <= 16'h803e;
		    ms <= ms_14;
		end
		ms_14: begin
		    q <= 16'h8043;
		    ms <= ms_15;
		end
		ms_15: begin
		    q <= 16'h8048;
		    ms <= ms_16;
		end
		ms_16: begin
		    q <= 16'h804d;
		    ms <= ms_17;
		end
		ms_17: begin
		    q <= 16'h8052;
		    ms <= ms_18;
		end
		ms_18: begin
		    q <= 16'h8057;
		    ms <= ms_19;
		end
		ms_19: begin
		    q <= 16'h805c;
		    ms <= ms_20;
		end
		ms_20: begin
		    q <= 16'h8061;
		    ms <= ms_21;
		end
		ms_21: begin
		    q <= 16'h8067;
		    ms <= ms_22;
		end
		ms_22: begin
		    q <= 16'h806c;
		    ms <= ms_23;
		end
		ms_23: begin
		    q <= 16'h8071;
		    ms <= ms_24;
		end
		ms_24: begin
		    q <= 16'h8076;
		    ms <= ms_25;
		end
		ms_25: begin
		    q <= 16'h807b;
		    ms <= ms_26;
		end
		ms_26: begin
		    q <= 16'h8080;
		    ms <= ms_27;
		end
		ms_27: begin
		    q <= 16'h8085;
		    ms <= ms_28;
		end
		ms_28: begin
		    q <= 16'h808a;
		    ms <= ms_29;
		end
		ms_29: begin
		    q <= 16'h808f;
		    ms <= ms_30;
		end
		ms_30: begin
		    q <= 16'h8094;
		    ms <= ms_31;
		end
		ms_31: begin
		    q <= 16'h8099;
		    ms <= ms_32;
		end
		ms_32: begin
		    q <= 16'h809e;
		    ms <= ms_33;
		end
		ms_33: begin
		    q <= 16'h80a3;
		    ms <= ms_34;
		end
		ms_34: begin
		    q <= 16'h80a8;
		    ms <= ms_35;
		end
		ms_35: begin
		    q <= 16'h80ad;
		    ms <= ms_36;
		end
		ms_36: begin
		    q <= 16'h80b2;
		    ms <= ms_37;
		end
		ms_37: begin
		    q <= 16'h80b7;
		    ms <= ms_38;
		end
		ms_38: begin
		    q <= 16'h80bc;
		    ms <= ms_39;
		end
		ms_39: begin
		    q <= 16'h80c1;
		    ms <= ms_40;
		end
		ms_40: begin
		    q <= 16'h80c6;
		    ms <= ms_41;
		end
		ms_41: begin
		    q <= 16'h80cb;
		    ms <= ms_42;
		end
		ms_42: begin
		    q <= 16'h80cf;
		    ms <= ms_43;
		end
		ms_43: begin
		    q <= 16'h80d4;
		    ms <= ms_44;
		end
		ms_44: begin
		    q <= 16'h80d9;
		    ms <= ms_45;
		end
		ms_45: begin
		    q <= 16'h80de;
		    ms <= ms_46;
		end
		ms_46: begin
		    q <= 16'h80e3;
		    ms <= ms_47;
		end
		ms_47: begin
		    q <= 16'h80e8;
		    ms <= ms_48;
		end
		ms_48: begin
		    q <= 16'h80ec;
		    ms <= ms_49;
		end
		ms_49: begin
		    q <= 16'h80f1;
		    ms <= ms_50;
		end
		ms_50: begin
		    q <= 16'h80f6;
		    ms <= ms_51;
		end
		ms_51: begin
		    q <= 16'h80fb;
		    ms <= ms_52;
		end
		ms_52: begin
		    q <= 16'h8100;
		    ms <= ms_53;
		end
		ms_53: begin
		    q <= 16'h8104;
		    ms <= ms_54;
		end
		ms_54: begin
		    q <= 16'h8109;
		    ms <= ms_55;
		end
		ms_55: begin
		    q <= 16'h810e;
		    ms <= ms_56;
		end
		ms_56: begin
		    q <= 16'h8112;
		    ms <= ms_57;
		end
		ms_57: begin
		    q <= 16'h8117;
		    ms <= ms_58;
		end
		ms_58: begin
		    q <= 16'h811c;
		    ms <= ms_59;
		end
		ms_59: begin
		    q <= 16'h8120;
		    ms <= ms_60;
		end
		ms_60: begin
		    q <= 16'h8125;
		    ms <= ms_61;
		end
		ms_61: begin
		    q <= 16'h812a;
		    ms <= ms_62;
		end
		ms_62: begin
		    q <= 16'h812e;
		    ms <= ms_63;
		end
		ms_63: begin
		    q <= 16'h8133;
		    ms <= ms_64;
		end
		ms_64: begin
		    q <= 16'h8137;
		    ms <= ms_65;
		end
		ms_65: begin
		    q <= 16'h813c;
		    ms <= ms_66;
		end
		ms_66: begin
		    q <= 16'h8140;
		    ms <= ms_67;
		end
		ms_67: begin
		    q <= 16'h8145;
		    ms <= ms_68;
		end
		ms_68: begin
		    q <= 16'h8149;
		    ms <= ms_69;
		end
		ms_69: begin
		    q <= 16'h814e;
		    ms <= ms_70;
		end
		ms_70: begin
		    q <= 16'h8152;
		    ms <= ms_71;
		end
		ms_71: begin
		    q <= 16'h8156;
		    ms <= ms_72;
		end
		ms_72: begin
		    q <= 16'h815b;
		    ms <= ms_73;
		end
		ms_73: begin
		    q <= 16'h815f;
		    ms <= ms_74;
		end
		ms_74: begin
		    q <= 16'h8163;
		    ms <= ms_75;
		end
		ms_75: begin
		    q <= 16'h8168;
		    ms <= ms_76;
		end
		ms_76: begin
		    q <= 16'h816c;
		    ms <= ms_77;
		end
		ms_77: begin
		    q <= 16'h8170;
		    ms <= ms_78;
		end
		ms_78: begin
		    q <= 16'h8175;
		    ms <= ms_79;
		end
		ms_79: begin
		    q <= 16'h8179;
		    ms <= ms_80;
		end
		ms_80: begin
		    q <= 16'h817d;
		    ms <= ms_81;
		end
		ms_81: begin
		    q <= 16'h8181;
		    ms <= ms_82;
		end
		ms_82: begin
		    q <= 16'h8185;
		    ms <= ms_83;
		end
		ms_83: begin
		    q <= 16'h8189;
		    ms <= ms_84;
		end
		ms_84: begin
		    q <= 16'h818e;
		    ms <= ms_85;
		end
		ms_85: begin
		    q <= 16'h8192;
		    ms <= ms_86;
		end
		ms_86: begin
		    q <= 16'h8196;
		    ms <= ms_87;
		end
		ms_87: begin
		    q <= 16'h819a;
		    ms <= ms_88;
		end
		ms_88: begin
		    q <= 16'h819e;
		    ms <= ms_89;
		end
		ms_89: begin
		    q <= 16'h81a2;
		    ms <= ms_90;
		end
		ms_90: begin
		    q <= 16'h81a6;
		    ms <= ms_91;
		end
		ms_91: begin
		    q <= 16'h81aa;
		    ms <= ms_92;
		end
		ms_92: begin
		    q <= 16'h81ae;
		    ms <= ms_93;
		end
		ms_93: begin
		    q <= 16'h81b1;
		    ms <= ms_94;
		end
		ms_94: begin
		    q <= 16'h81b5;
		    ms <= ms_95;
		end
		ms_95: begin
		    q <= 16'h81b9;
		    ms <= ms_96;
		end
		ms_96: begin
		    q <= 16'h81bd;
		    ms <= ms_97;
		end
		ms_97: begin
		    q <= 16'h81c1;
		    ms <= ms_98;
		end
		ms_98: begin
		    q <= 16'h81c4;
		    ms <= ms_99;
		end
		ms_99: begin
		    q <= 16'h81c8;
		    ms <= ms_100;
		end
		ms_100: begin
		    q <= 16'h81cc;
		    ms <= ms_101;
		end
		ms_101: begin
		    q <= 16'h81cf;
		    ms <= ms_102;
		end
		ms_102: begin
		    q <= 16'h81d3;
		    ms <= ms_103;
		end
		ms_103: begin
		    q <= 16'h81d7;
		    ms <= ms_104;
		end
		ms_104: begin
		    q <= 16'h81da;
		    ms <= ms_105;
		end
		ms_105: begin
		    q <= 16'h81de;
		    ms <= ms_106;
		end
		ms_106: begin
		    q <= 16'h81e1;
		    ms <= ms_107;
		end
		ms_107: begin
		    q <= 16'h81e5;
		    ms <= ms_108;
		end
		ms_108: begin
		    q <= 16'h81e8;
		    ms <= ms_109;
		end
		ms_109: begin
		    q <= 16'h81ec;
		    ms <= ms_110;
		end
		ms_110: begin
		    q <= 16'h81ef;
		    ms <= ms_111;
		end
		ms_111: begin
		    q <= 16'h81f2;
		    ms <= ms_112;
		end
		ms_112: begin
		    q <= 16'h81f6;
		    ms <= ms_113;
		end
		ms_113: begin
		    q <= 16'h81f9;
		    ms <= ms_114;
		end
		ms_114: begin
		    q <= 16'h81fc;
		    ms <= ms_115;
		end
		ms_115: begin
		    q <= 16'h81ff;
		    ms <= ms_116;
		end
		ms_116: begin
		    q <= 16'h8203;
		    ms <= ms_117;
		end
		ms_117: begin
		    q <= 16'h8206;
		    ms <= ms_118;
		end
		ms_118: begin
		    q <= 16'h8209;
		    ms <= ms_119;
		end
		ms_119: begin
		    q <= 16'h820c;
		    ms <= ms_120;
		end
		ms_120: begin
		    q <= 16'h820f;
		    ms <= ms_121;
		end
		ms_121: begin
		    q <= 16'h8212;
		    ms <= ms_122;
		end
		ms_122: begin
		    q <= 16'h8215;
		    ms <= ms_123;
		end
		ms_123: begin
		    q <= 16'h8218;
		    ms <= ms_124;
		end
		ms_124: begin
		    q <= 16'h821b;
		    ms <= ms_125;
		end
		ms_125: begin
		    q <= 16'h821e;
		    ms <= ms_126;
		end
		ms_126: begin
		    q <= 16'h8221;
		    ms <= ms_127;
		end
		ms_127: begin
		    q <= 16'h8224;
		    ms <= ms_128;
		end
		ms_128: begin
		    q <= 16'h8227;
		    ms <= ms_129;
		end
		ms_129: begin
		    q <= 16'h8229;
		    ms <= ms_130;
		end
		ms_130: begin
		    q <= 16'h822c;
		    ms <= ms_131;
		end
		ms_131: begin
		    q <= 16'h822f;
		    ms <= ms_132;
		end
		ms_132: begin
		    q <= 16'h8231;
		    ms <= ms_133;
		end
		ms_133: begin
		    q <= 16'h8234;
		    ms <= ms_134;
		end
		ms_134: begin
		    q <= 16'h8237;
		    ms <= ms_135;
		end
		ms_135: begin
		    q <= 16'h8239;
		    ms <= ms_136;
		end
		ms_136: begin
		    q <= 16'h823c;
		    ms <= ms_137;
		end
		ms_137: begin
		    q <= 16'h823e;
		    ms <= ms_138;
		end
		ms_138: begin
		    q <= 16'h8241;
		    ms <= ms_139;
		end
		ms_139: begin
		    q <= 16'h8243;
		    ms <= ms_140;
		end
		ms_140: begin
		    q <= 16'h8246;
		    ms <= ms_141;
		end
		ms_141: begin
		    q <= 16'h8248;
		    ms <= ms_142;
		end
		ms_142: begin
		    q <= 16'h824a;
		    ms <= ms_143;
		end
		ms_143: begin
		    q <= 16'h824d;
		    ms <= ms_144;
		end
		ms_144: begin
		    q <= 16'h824f;
		    ms <= ms_145;
		end
		ms_145: begin
		    q <= 16'h8251;
		    ms <= ms_146;
		end
		ms_146: begin
		    q <= 16'h8253;
		    ms <= ms_147;
		end
		ms_147: begin
		    q <= 16'h8255;
		    ms <= ms_148;
		end
		ms_148: begin
		    q <= 16'h8257;
		    ms <= ms_149;
		end
		ms_149: begin
		    q <= 16'h8259;
		    ms <= ms_150;
		end
		ms_150: begin
		    q <= 16'h825b;
		    ms <= ms_151;
		end
		ms_151: begin
		    q <= 16'h825d;
		    ms <= ms_152;
		end
		ms_152: begin
		    q <= 16'h825f;
		    ms <= ms_153;
		end
		ms_153: begin
		    q <= 16'h8261;
		    ms <= ms_154;
		end
		ms_154: begin
		    q <= 16'h8263;
		    ms <= ms_155;
		end
		ms_155: begin
		    q <= 16'h8265;
		    ms <= ms_156;
		end
		ms_156: begin
		    q <= 16'h8267;
		    ms <= ms_157;
		end
		ms_157: begin
		    q <= 16'h8269;
		    ms <= ms_158;
		end
		ms_158: begin
		    q <= 16'h826a;
		    ms <= ms_159;
		end
		ms_159: begin
		    q <= 16'h826c;
		    ms <= ms_160;
		end
		ms_160: begin
		    q <= 16'h826e;
		    ms <= ms_161;
		end
		ms_161: begin
		    q <= 16'h826f;
		    ms <= ms_162;
		end
		ms_162: begin
		    q <= 16'h8271;
		    ms <= ms_163;
		end
		ms_163: begin
		    q <= 16'h8272;
		    ms <= ms_164;
		end
		ms_164: begin
		    q <= 16'h8274;
		    ms <= ms_165;
		end
		ms_165: begin
		    q <= 16'h8275;
		    ms <= ms_166;
		end
		ms_166: begin
		    q <= 16'h8277;
		    ms <= ms_167;
		end
		ms_167: begin
		    q <= 16'h8278;
		    ms <= ms_168;
		end
		ms_168: begin
		    q <= 16'h8279;
		    ms <= ms_169;
		end
		ms_169: begin
		    q <= 16'h827b;
		    ms <= ms_170;
		end
		ms_170: begin
		    q <= 16'h827c;
		    ms <= ms_171;
		end
		ms_171: begin
		    q <= 16'h827d;
		    ms <= ms_172;
		end
		ms_172: begin
		    q <= 16'h827e;
		    ms <= ms_173;
		end
		ms_173: begin
		    q <= 16'h8280;
		    ms <= ms_174;
		end
		ms_174: begin
		    q <= 16'h8281;
		    ms <= ms_175;
		end
		ms_175: begin
		    q <= 16'h8282;
		    ms <= ms_176;
		end
		ms_176: begin
		    q <= 16'h8283;
		    ms <= ms_177;
		end
		ms_177: begin
		    q <= 16'h8284;
		    ms <= ms_178;
		end
		ms_178: begin
		    q <= 16'h8285;
		    ms <= ms_179;
		end
		ms_179: begin
		    q <= 16'h8286;
		    ms <= ms_180;
		end
		ms_180: begin
		    q <= 16'h8286;
		    ms <= ms_181;
		end
		ms_181: begin
		    q <= 16'h8287;
		    ms <= ms_182;
		end
		ms_182: begin
		    q <= 16'h8288;
		    ms <= ms_183;
		end
		ms_183: begin
		    q <= 16'h8289;
		    ms <= ms_184;
		end
		ms_184: begin
		    q <= 16'h828a;
		    ms <= ms_185;
		end
		ms_185: begin
		    q <= 16'h828a;
		    ms <= ms_186;
		end
		ms_186: begin
		    q <= 16'h828b;
		    ms <= ms_187;
		end
		ms_187: begin
		    q <= 16'h828b;
		    ms <= ms_188;
		end
		ms_188: begin
		    q <= 16'h828c;
		    ms <= ms_189;
		end
		ms_189: begin
		    q <= 16'h828c;
		    ms <= ms_190;
		end
		ms_190: begin
		    q <= 16'h828d;
		    ms <= ms_191;
		end
		ms_191: begin
		    q <= 16'h828d;
		    ms <= ms_192;
		end
		ms_192: begin
		    q <= 16'h828e;
		    ms <= ms_193;
		end
		ms_193: begin
		    q <= 16'h828e;
		    ms <= ms_194;
		end
		ms_194: begin
		    q <= 16'h828e;
		    ms <= ms_195;
		end
		ms_195: begin
		    q <= 16'h828f;
		    ms <= ms_196;
		end
		ms_196: begin
		    q <= 16'h828f;
		    ms <= ms_197;
		end
		ms_197: begin
		    q <= 16'h828f;
		    ms <= ms_198;
		end
		ms_198: begin
		    q <= 16'h828f;
		    ms <= ms_199;
		end
		ms_199: begin
		    q <= 16'h828f;
		    ms <= ms_200;
		end
		ms_200: begin
		    q <= 16'h828f;
		    ms <= ms_201;
		end
		ms_201: begin
		    q <= 16'h828f;
		    ms <= ms_202;
		end
		ms_202: begin
		    q <= 16'h828f;
		    ms <= ms_203;
		end
		ms_203: begin
		    q <= 16'h828f;
		    ms <= ms_204;
		end
		ms_204: begin
		    q <= 16'h828f;
		    ms <= ms_205;
		end
		ms_205: begin
		    q <= 16'h828f;
		    ms <= ms_206;
		end
		ms_206: begin
		    q <= 16'h828f;
		    ms <= ms_207;
		end
		ms_207: begin
		    q <= 16'h828f;
		    ms <= ms_208;
		end
		ms_208: begin
		    q <= 16'h828e;
		    ms <= ms_209;
		end
		ms_209: begin
		    q <= 16'h828e;
		    ms <= ms_210;
		end
		ms_210: begin
		    q <= 16'h828e;
		    ms <= ms_211;
		end
		ms_211: begin
		    q <= 16'h828d;
		    ms <= ms_212;
		end
		ms_212: begin
		    q <= 16'h828d;
		    ms <= ms_213;
		end
		ms_213: begin
		    q <= 16'h828c;
		    ms <= ms_214;
		end
		ms_214: begin
		    q <= 16'h828c;
		    ms <= ms_215;
		end
		ms_215: begin
		    q <= 16'h828b;
		    ms <= ms_216;
		end
		ms_216: begin
		    q <= 16'h828b;
		    ms <= ms_217;
		end
		ms_217: begin
		    q <= 16'h828a;
		    ms <= ms_218;
		end
		ms_218: begin
		    q <= 16'h828a;
		    ms <= ms_219;
		end
		ms_219: begin
		    q <= 16'h8289;
		    ms <= ms_220;
		end
		ms_220: begin
		    q <= 16'h8288;
		    ms <= ms_221;
		end
		ms_221: begin
		    q <= 16'h8287;
		    ms <= ms_222;
		end
		ms_222: begin
		    q <= 16'h8286;
		    ms <= ms_223;
		end
		ms_223: begin
		    q <= 16'h8286;
		    ms <= ms_224;
		end
		ms_224: begin
		    q <= 16'h8285;
		    ms <= ms_225;
		end
		ms_225: begin
		    q <= 16'h8284;
		    ms <= ms_226;
		end
		ms_226: begin
		    q <= 16'h8283;
		    ms <= ms_227;
		end
		ms_227: begin
		    q <= 16'h8282;
		    ms <= ms_228;
		end
		ms_228: begin
		    q <= 16'h8281;
		    ms <= ms_229;
		end
		ms_229: begin
		    q <= 16'h8280;
		    ms <= ms_230;
		end
		ms_230: begin
		    q <= 16'h827e;
		    ms <= ms_231;
		end
		ms_231: begin
		    q <= 16'h827d;
		    ms <= ms_232;
		end
		ms_232: begin
		    q <= 16'h827c;
		    ms <= ms_233;
		end
		ms_233: begin
		    q <= 16'h827b;
		    ms <= ms_234;
		end
		ms_234: begin
		    q <= 16'h8279;
		    ms <= ms_235;
		end
		ms_235: begin
		    q <= 16'h8278;
		    ms <= ms_236;
		end
		ms_236: begin
		    q <= 16'h8277;
		    ms <= ms_237;
		end
		ms_237: begin
		    q <= 16'h8275;
		    ms <= ms_238;
		end
		ms_238: begin
		    q <= 16'h8274;
		    ms <= ms_239;
		end
		ms_239: begin
		    q <= 16'h8272;
		    ms <= ms_240;
		end
		ms_240: begin
		    q <= 16'h8271;
		    ms <= ms_241;
		end
		ms_241: begin
		    q <= 16'h826f;
		    ms <= ms_242;
		end
		ms_242: begin
		    q <= 16'h826e;
		    ms <= ms_243;
		end
		ms_243: begin
		    q <= 16'h826c;
		    ms <= ms_244;
		end
		ms_244: begin
		    q <= 16'h826a;
		    ms <= ms_245;
		end
		ms_245: begin
		    q <= 16'h8269;
		    ms <= ms_246;
		end
		ms_246: begin
		    q <= 16'h8267;
		    ms <= ms_247;
		end
		ms_247: begin
		    q <= 16'h8265;
		    ms <= ms_248;
		end
		ms_248: begin
		    q <= 16'h8263;
		    ms <= ms_249;
		end
		ms_249: begin
		    q <= 16'h8261;
		    ms <= ms_250;
		end
		ms_250: begin
		    q <= 16'h825f;
		    ms <= ms_251;
		end
		ms_251: begin
		    q <= 16'h825d;
		    ms <= ms_252;
		end
		ms_252: begin
		    q <= 16'h825b;
		    ms <= ms_253;
		end
		ms_253: begin
		    q <= 16'h8259;
		    ms <= ms_254;
		end
		ms_254: begin
		    q <= 16'h8257;
		    ms <= ms_255;
		end
		ms_255: begin
		    q <= 16'h8255;
		    ms <= ms_256;
		end
		ms_256: begin
		    q <= 16'h8253;
		    ms <= ms_257;
		end
		ms_257: begin
		    q <= 16'h8251;
		    ms <= ms_258;
		end
		ms_258: begin
		    q <= 16'h824f;
		    ms <= ms_259;
		end
		ms_259: begin
		    q <= 16'h824d;
		    ms <= ms_260;
		end
		ms_260: begin
		    q <= 16'h824a;
		    ms <= ms_261;
		end
		ms_261: begin
		    q <= 16'h8248;
		    ms <= ms_262;
		end
		ms_262: begin
		    q <= 16'h8246;
		    ms <= ms_263;
		end
		ms_263: begin
		    q <= 16'h8243;
		    ms <= ms_264;
		end
		ms_264: begin
		    q <= 16'h8241;
		    ms <= ms_265;
		end
		ms_265: begin
		    q <= 16'h823e;
		    ms <= ms_266;
		end
		ms_266: begin
		    q <= 16'h823c;
		    ms <= ms_267;
		end
		ms_267: begin
		    q <= 16'h8239;
		    ms <= ms_268;
		end
		ms_268: begin
		    q <= 16'h8237;
		    ms <= ms_269;
		end
		ms_269: begin
		    q <= 16'h8234;
		    ms <= ms_270;
		end
		ms_270: begin
		    q <= 16'h8231;
		    ms <= ms_271;
		end
		ms_271: begin
		    q <= 16'h822f;
		    ms <= ms_272;
		end
		ms_272: begin
		    q <= 16'h822c;
		    ms <= ms_273;
		end
		ms_273: begin
		    q <= 16'h8229;
		    ms <= ms_274;
		end
		ms_274: begin
		    q <= 16'h8227;
		    ms <= ms_275;
		end
		ms_275: begin
		    q <= 16'h8224;
		    ms <= ms_276;
		end
		ms_276: begin
		    q <= 16'h8221;
		    ms <= ms_277;
		end
		ms_277: begin
		    q <= 16'h821e;
		    ms <= ms_278;
		end
		ms_278: begin
		    q <= 16'h821b;
		    ms <= ms_279;
		end
		ms_279: begin
		    q <= 16'h8218;
		    ms <= ms_280;
		end
		ms_280: begin
		    q <= 16'h8215;
		    ms <= ms_281;
		end
		ms_281: begin
		    q <= 16'h8212;
		    ms <= ms_282;
		end
		ms_282: begin
		    q <= 16'h820f;
		    ms <= ms_283;
		end
		ms_283: begin
		    q <= 16'h820c;
		    ms <= ms_284;
		end
		ms_284: begin
		    q <= 16'h8209;
		    ms <= ms_285;
		end
		ms_285: begin
		    q <= 16'h8206;
		    ms <= ms_286;
		end
		ms_286: begin
		    q <= 16'h8203;
		    ms <= ms_287;
		end
		ms_287: begin
		    q <= 16'h81ff;
		    ms <= ms_288;
		end
		ms_288: begin
		    q <= 16'h81fc;
		    ms <= ms_289;
		end
		ms_289: begin
		    q <= 16'h81f9;
		    ms <= ms_290;
		end
		ms_290: begin
		    q <= 16'h81f6;
		    ms <= ms_291;
		end
		ms_291: begin
		    q <= 16'h81f2;
		    ms <= ms_292;
		end
		ms_292: begin
		    q <= 16'h81ef;
		    ms <= ms_293;
		end
		ms_293: begin
		    q <= 16'h81ec;
		    ms <= ms_294;
		end
		ms_294: begin
		    q <= 16'h81e8;
		    ms <= ms_295;
		end
		ms_295: begin
		    q <= 16'h81e5;
		    ms <= ms_296;
		end
		ms_296: begin
		    q <= 16'h81e1;
		    ms <= ms_297;
		end
		ms_297: begin
		    q <= 16'h81de;
		    ms <= ms_298;
		end
		ms_298: begin
		    q <= 16'h81da;
		    ms <= ms_299;
		end
		ms_299: begin
		    q <= 16'h81d7;
		    ms <= ms_300;
		end
		ms_300: begin
		    q <= 16'h81d3;
		    ms <= ms_301;
		end
		ms_301: begin
		    q <= 16'h81cf;
		    ms <= ms_302;
		end
		ms_302: begin
		    q <= 16'h81cc;
		    ms <= ms_303;
		end
		ms_303: begin
		    q <= 16'h81c8;
		    ms <= ms_304;
		end
		ms_304: begin
		    q <= 16'h81c4;
		    ms <= ms_305;
		end
		ms_305: begin
		    q <= 16'h81c1;
		    ms <= ms_306;
		end
		ms_306: begin
		    q <= 16'h81bd;
		    ms <= ms_307;
		end
		ms_307: begin
		    q <= 16'h81b9;
		    ms <= ms_308;
		end
		ms_308: begin
		    q <= 16'h81b5;
		    ms <= ms_309;
		end
		ms_309: begin
		    q <= 16'h81b1;
		    ms <= ms_310;
		end
		ms_310: begin
		    q <= 16'h81ae;
		    ms <= ms_311;
		end
		ms_311: begin
		    q <= 16'h81aa;
		    ms <= ms_312;
		end
		ms_312: begin
		    q <= 16'h81a6;
		    ms <= ms_313;
		end
		ms_313: begin
		    q <= 16'h81a2;
		    ms <= ms_314;
		end
		ms_314: begin
		    q <= 16'h819e;
		    ms <= ms_315;
		end
		ms_315: begin
		    q <= 16'h819a;
		    ms <= ms_316;
		end
		ms_316: begin
		    q <= 16'h8196;
		    ms <= ms_317;
		end
		ms_317: begin
		    q <= 16'h8192;
		    ms <= ms_318;
		end
		ms_318: begin
		    q <= 16'h818e;
		    ms <= ms_319;
		end
		ms_319: begin
		    q <= 16'h8189;
		    ms <= ms_320;
		end
		ms_320: begin
		    q <= 16'h8185;
		    ms <= ms_321;
		end
		ms_321: begin
		    q <= 16'h8181;
		    ms <= ms_322;
		end
		ms_322: begin
		    q <= 16'h817d;
		    ms <= ms_323;
		end
		ms_323: begin
		    q <= 16'h8179;
		    ms <= ms_324;
		end
		ms_324: begin
		    q <= 16'h8175;
		    ms <= ms_325;
		end
		ms_325: begin
		    q <= 16'h8170;
		    ms <= ms_326;
		end
		ms_326: begin
		    q <= 16'h816c;
		    ms <= ms_327;
		end
		ms_327: begin
		    q <= 16'h8168;
		    ms <= ms_328;
		end
		ms_328: begin
		    q <= 16'h8163;
		    ms <= ms_329;
		end
		ms_329: begin
		    q <= 16'h815f;
		    ms <= ms_330;
		end
		ms_330: begin
		    q <= 16'h815b;
		    ms <= ms_331;
		end
		ms_331: begin
		    q <= 16'h8156;
		    ms <= ms_332;
		end
		ms_332: begin
		    q <= 16'h8152;
		    ms <= ms_333;
		end
		ms_333: begin
		    q <= 16'h814e;
		    ms <= ms_334;
		end
		ms_334: begin
		    q <= 16'h8149;
		    ms <= ms_335;
		end
		ms_335: begin
		    q <= 16'h8145;
		    ms <= ms_336;
		end
		ms_336: begin
		    q <= 16'h8140;
		    ms <= ms_337;
		end
		ms_337: begin
		    q <= 16'h813c;
		    ms <= ms_338;
		end
		ms_338: begin
		    q <= 16'h8137;
		    ms <= ms_339;
		end
		ms_339: begin
		    q <= 16'h8133;
		    ms <= ms_340;
		end
		ms_340: begin
		    q <= 16'h812e;
		    ms <= ms_341;
		end
		ms_341: begin
		    q <= 16'h812a;
		    ms <= ms_342;
		end
		ms_342: begin
		    q <= 16'h8125;
		    ms <= ms_343;
		end
		ms_343: begin
		    q <= 16'h8120;
		    ms <= ms_344;
		end
		ms_344: begin
		    q <= 16'h811c;
		    ms <= ms_345;
		end
		ms_345: begin
		    q <= 16'h8117;
		    ms <= ms_346;
		end
		ms_346: begin
		    q <= 16'h8112;
		    ms <= ms_347;
		end
		ms_347: begin
		    q <= 16'h810e;
		    ms <= ms_348;
		end
		ms_348: begin
		    q <= 16'h8109;
		    ms <= ms_349;
		end
		ms_349: begin
		    q <= 16'h8104;
		    ms <= ms_350;
		end
		ms_350: begin
		    q <= 16'h8100;
		    ms <= ms_351;
		end
		ms_351: begin
		    q <= 16'h80fb;
		    ms <= ms_352;
		end
		ms_352: begin
		    q <= 16'h80f6;
		    ms <= ms_353;
		end
		ms_353: begin
		    q <= 16'h80f1;
		    ms <= ms_354;
		end
		ms_354: begin
		    q <= 16'h80ec;
		    ms <= ms_355;
		end
		ms_355: begin
		    q <= 16'h80e8;
		    ms <= ms_356;
		end
		ms_356: begin
		    q <= 16'h80e3;
		    ms <= ms_357;
		end
		ms_357: begin
		    q <= 16'h80de;
		    ms <= ms_358;
		end
		ms_358: begin
		    q <= 16'h80d9;
		    ms <= ms_359;
		end
		ms_359: begin
		    q <= 16'h80d4;
		    ms <= ms_360;
		end
		ms_360: begin
		    q <= 16'h80cf;
		    ms <= ms_361;
		end
		ms_361: begin
		    q <= 16'h80cb;
		    ms <= ms_362;
		end
		ms_362: begin
		    q <= 16'h80c6;
		    ms <= ms_363;
		end
		ms_363: begin
		    q <= 16'h80c1;
		    ms <= ms_364;
		end
		ms_364: begin
		    q <= 16'h80bc;
		    ms <= ms_365;
		end
		ms_365: begin
		    q <= 16'h80b7;
		    ms <= ms_366;
		end
		ms_366: begin
		    q <= 16'h80b2;
		    ms <= ms_367;
		end
		ms_367: begin
		    q <= 16'h80ad;
		    ms <= ms_368;
		end
		ms_368: begin
		    q <= 16'h80a8;
		    ms <= ms_369;
		end
		ms_369: begin
		    q <= 16'h80a3;
		    ms <= ms_370;
		end
		ms_370: begin
		    q <= 16'h809e;
		    ms <= ms_371;
		end
		ms_371: begin
		    q <= 16'h8099;
		    ms <= ms_372;
		end
		ms_372: begin
		    q <= 16'h8094;
		    ms <= ms_373;
		end
		ms_373: begin
		    q <= 16'h808f;
		    ms <= ms_374;
		end
		ms_374: begin
		    q <= 16'h808a;
		    ms <= ms_375;
		end
		ms_375: begin
		    q <= 16'h8085;
		    ms <= ms_376;
		end
		ms_376: begin
		    q <= 16'h8080;
		    ms <= ms_377;
		end
		ms_377: begin
		    q <= 16'h807b;
		    ms <= ms_378;
		end
		ms_378: begin
		    q <= 16'h8076;
		    ms <= ms_379;
		end
		ms_379: begin
		    q <= 16'h8071;
		    ms <= ms_380;
		end
		ms_380: begin
		    q <= 16'h806c;
		    ms <= ms_381;
		end
		ms_381: begin
		    q <= 16'h8067;
		    ms <= ms_382;
		end
		ms_382: begin
		    q <= 16'h8061;
		    ms <= ms_383;
		end
		ms_383: begin
		    q <= 16'h805c;
		    ms <= ms_384;
		end
		ms_384: begin
		    q <= 16'h8057;
		    ms <= ms_385;
		end
		ms_385: begin
		    q <= 16'h8052;
		    ms <= ms_386;
		end
		ms_386: begin
		    q <= 16'h804d;
		    ms <= ms_387;
		end
		ms_387: begin
		    q <= 16'h8048;
		    ms <= ms_388;
		end
		ms_388: begin
		    q <= 16'h8043;
		    ms <= ms_389;
		end
		ms_389: begin
		    q <= 16'h803e;
		    ms <= ms_390;
		end
		ms_390: begin
		    q <= 16'h8039;
		    ms <= ms_391;
		end
		ms_391: begin
		    q <= 16'h8033;
		    ms <= ms_392;
		end
		ms_392: begin
		    q <= 16'h802e;
		    ms <= ms_393;
		end
		ms_393: begin
		    q <= 16'h8029;
		    ms <= ms_394;
		end
		ms_394: begin
		    q <= 16'h8024;
		    ms <= ms_395;
		end
		ms_395: begin
		    q <= 16'h801f;
		    ms <= ms_396;
		end
		ms_396: begin
		    q <= 16'h801a;
		    ms <= ms_397;
		end
		ms_397: begin
		    q <= 16'h8015;
		    ms <= ms_398;
		end
		ms_398: begin
		    q <= 16'h800f;
		    ms <= ms_399;
		end
		ms_399: begin
		    q <= 16'h800a;
		    ms <= ms_400;
		end
		ms_400: begin
		    q <= 16'h8005;
		    ms <= ms_401;
		end
		ms_401: begin
		    q <= 16'h8000;
		    ms <= ms_402;
		end
		ms_402: begin
		    q <= 16'h7ffb;
		    ms <= ms_403;
		end
		ms_403: begin
		    q <= 16'h7ff6;
		    ms <= ms_404;
		end
		ms_404: begin
		    q <= 16'h7ff1;
		    ms <= ms_405;
		end
		ms_405: begin
		    q <= 16'h7feb;
		    ms <= ms_406;
		end
		ms_406: begin
		    q <= 16'h7fe6;
		    ms <= ms_407;
		end
		ms_407: begin
		    q <= 16'h7fe1;
		    ms <= ms_408;
		end
		ms_408: begin
		    q <= 16'h7fdc;
		    ms <= ms_409;
		end
		ms_409: begin
		    q <= 16'h7fd7;
		    ms <= ms_410;
		end
		ms_410: begin
		    q <= 16'h7fd2;
		    ms <= ms_411;
		end
		ms_411: begin
		    q <= 16'h7fcd;
		    ms <= ms_412;
		end
		ms_412: begin
		    q <= 16'h7fc7;
		    ms <= ms_413;
		end
		ms_413: begin
		    q <= 16'h7fc2;
		    ms <= ms_414;
		end
		ms_414: begin
		    q <= 16'h7fbd;
		    ms <= ms_415;
		end
		ms_415: begin
		    q <= 16'h7fb8;
		    ms <= ms_416;
		end
		ms_416: begin
		    q <= 16'h7fb3;
		    ms <= ms_417;
		end
		ms_417: begin
		    q <= 16'h7fae;
		    ms <= ms_418;
		end
		ms_418: begin
		    q <= 16'h7fa9;
		    ms <= ms_419;
		end
		ms_419: begin
		    q <= 16'h7fa4;
		    ms <= ms_420;
		end
		ms_420: begin
		    q <= 16'h7f9f;
		    ms <= ms_421;
		end
		ms_421: begin
		    q <= 16'h7f99;
		    ms <= ms_422;
		end
		ms_422: begin
		    q <= 16'h7f94;
		    ms <= ms_423;
		end
		ms_423: begin
		    q <= 16'h7f8f;
		    ms <= ms_424;
		end
		ms_424: begin
		    q <= 16'h7f8a;
		    ms <= ms_425;
		end
		ms_425: begin
		    q <= 16'h7f85;
		    ms <= ms_426;
		end
		ms_426: begin
		    q <= 16'h7f80;
		    ms <= ms_427;
		end
		ms_427: begin
		    q <= 16'h7f7b;
		    ms <= ms_428;
		end
		ms_428: begin
		    q <= 16'h7f76;
		    ms <= ms_429;
		end
		ms_429: begin
		    q <= 16'h7f71;
		    ms <= ms_430;
		end
		ms_430: begin
		    q <= 16'h7f6c;
		    ms <= ms_431;
		end
		ms_431: begin
		    q <= 16'h7f67;
		    ms <= ms_432;
		end
		ms_432: begin
		    q <= 16'h7f62;
		    ms <= ms_433;
		end
		ms_433: begin
		    q <= 16'h7f5d;
		    ms <= ms_434;
		end
		ms_434: begin
		    q <= 16'h7f58;
		    ms <= ms_435;
		end
		ms_435: begin
		    q <= 16'h7f53;
		    ms <= ms_436;
		end
		ms_436: begin
		    q <= 16'h7f4e;
		    ms <= ms_437;
		end
		ms_437: begin
		    q <= 16'h7f49;
		    ms <= ms_438;
		end
		ms_438: begin
		    q <= 16'h7f44;
		    ms <= ms_439;
		end
		ms_439: begin
		    q <= 16'h7f3f;
		    ms <= ms_440;
		end
		ms_440: begin
		    q <= 16'h7f3a;
		    ms <= ms_441;
		end
		ms_441: begin
		    q <= 16'h7f35;
		    ms <= ms_442;
		end
		ms_442: begin
		    q <= 16'h7f31;
		    ms <= ms_443;
		end
		ms_443: begin
		    q <= 16'h7f2c;
		    ms <= ms_444;
		end
		ms_444: begin
		    q <= 16'h7f27;
		    ms <= ms_445;
		end
		ms_445: begin
		    q <= 16'h7f22;
		    ms <= ms_446;
		end
		ms_446: begin
		    q <= 16'h7f1d;
		    ms <= ms_447;
		end
		ms_447: begin
		    q <= 16'h7f18;
		    ms <= ms_448;
		end
		ms_448: begin
		    q <= 16'h7f14;
		    ms <= ms_449;
		end
		ms_449: begin
		    q <= 16'h7f0f;
		    ms <= ms_450;
		end
		ms_450: begin
		    q <= 16'h7f0a;
		    ms <= ms_451;
		end
		ms_451: begin
		    q <= 16'h7f05;
		    ms <= ms_452;
		end
		ms_452: begin
		    q <= 16'h7f00;
		    ms <= ms_453;
		end
		ms_453: begin
		    q <= 16'h7efc;
		    ms <= ms_454;
		end
		ms_454: begin
		    q <= 16'h7ef7;
		    ms <= ms_455;
		end
		ms_455: begin
		    q <= 16'h7ef2;
		    ms <= ms_456;
		end
		ms_456: begin
		    q <= 16'h7eee;
		    ms <= ms_457;
		end
		ms_457: begin
		    q <= 16'h7ee9;
		    ms <= ms_458;
		end
		ms_458: begin
		    q <= 16'h7ee4;
		    ms <= ms_459;
		end
		ms_459: begin
		    q <= 16'h7ee0;
		    ms <= ms_460;
		end
		ms_460: begin
		    q <= 16'h7edb;
		    ms <= ms_461;
		end
		ms_461: begin
		    q <= 16'h7ed6;
		    ms <= ms_462;
		end
		ms_462: begin
		    q <= 16'h7ed2;
		    ms <= ms_463;
		end
		ms_463: begin
		    q <= 16'h7ecd;
		    ms <= ms_464;
		end
		ms_464: begin
		    q <= 16'h7ec9;
		    ms <= ms_465;
		end
		ms_465: begin
		    q <= 16'h7ec4;
		    ms <= ms_466;
		end
		ms_466: begin
		    q <= 16'h7ec0;
		    ms <= ms_467;
		end
		ms_467: begin
		    q <= 16'h7ebb;
		    ms <= ms_468;
		end
		ms_468: begin
		    q <= 16'h7eb7;
		    ms <= ms_469;
		end
		ms_469: begin
		    q <= 16'h7eb2;
		    ms <= ms_470;
		end
		ms_470: begin
		    q <= 16'h7eae;
		    ms <= ms_471;
		end
		ms_471: begin
		    q <= 16'h7eaa;
		    ms <= ms_472;
		end
		ms_472: begin
		    q <= 16'h7ea5;
		    ms <= ms_473;
		end
		ms_473: begin
		    q <= 16'h7ea1;
		    ms <= ms_474;
		end
		ms_474: begin
		    q <= 16'h7e9d;
		    ms <= ms_475;
		end
		ms_475: begin
		    q <= 16'h7e98;
		    ms <= ms_476;
		end
		ms_476: begin
		    q <= 16'h7e94;
		    ms <= ms_477;
		end
		ms_477: begin
		    q <= 16'h7e90;
		    ms <= ms_478;
		end
		ms_478: begin
		    q <= 16'h7e8b;
		    ms <= ms_479;
		end
		ms_479: begin
		    q <= 16'h7e87;
		    ms <= ms_480;
		end
		ms_480: begin
		    q <= 16'h7e83;
		    ms <= ms_481;
		end
		ms_481: begin
		    q <= 16'h7e7f;
		    ms <= ms_482;
		end
		ms_482: begin
		    q <= 16'h7e7b;
		    ms <= ms_483;
		end
		ms_483: begin
		    q <= 16'h7e77;
		    ms <= ms_484;
		end
		ms_484: begin
		    q <= 16'h7e72;
		    ms <= ms_485;
		end
		ms_485: begin
		    q <= 16'h7e6e;
		    ms <= ms_486;
		end
		ms_486: begin
		    q <= 16'h7e6a;
		    ms <= ms_487;
		end
		ms_487: begin
		    q <= 16'h7e66;
		    ms <= ms_488;
		end
		ms_488: begin
		    q <= 16'h7e62;
		    ms <= ms_489;
		end
		ms_489: begin
		    q <= 16'h7e5e;
		    ms <= ms_490;
		end
		ms_490: begin
		    q <= 16'h7e5a;
		    ms <= ms_491;
		end
		ms_491: begin
		    q <= 16'h7e56;
		    ms <= ms_492;
		end
		ms_492: begin
		    q <= 16'h7e52;
		    ms <= ms_493;
		end
		ms_493: begin
		    q <= 16'h7e4f;
		    ms <= ms_494;
		end
		ms_494: begin
		    q <= 16'h7e4b;
		    ms <= ms_495;
		end
		ms_495: begin
		    q <= 16'h7e47;
		    ms <= ms_496;
		end
		ms_496: begin
		    q <= 16'h7e43;
		    ms <= ms_497;
		end
		ms_497: begin
		    q <= 16'h7e3f;
		    ms <= ms_498;
		end
		ms_498: begin
		    q <= 16'h7e3c;
		    ms <= ms_499;
		end
		ms_499: begin
		    q <= 16'h7e38;
		    ms <= ms_500;
		end
		ms_500: begin
		    q <= 16'h7e34;
		    ms <= ms_501;
		end
		ms_501: begin
		    q <= 16'h7e31;
		    ms <= ms_502;
		end
		ms_502: begin
		    q <= 16'h7e2d;
		    ms <= ms_503;
		end
		ms_503: begin
		    q <= 16'h7e29;
		    ms <= ms_504;
		end
		ms_504: begin
		    q <= 16'h7e26;
		    ms <= ms_505;
		end
		ms_505: begin
		    q <= 16'h7e22;
		    ms <= ms_506;
		end
		ms_506: begin
		    q <= 16'h7e1f;
		    ms <= ms_507;
		end
		ms_507: begin
		    q <= 16'h7e1b;
		    ms <= ms_508;
		end
		ms_508: begin
		    q <= 16'h7e18;
		    ms <= ms_509;
		end
		ms_509: begin
		    q <= 16'h7e14;
		    ms <= ms_510;
		end
		ms_510: begin
		    q <= 16'h7e11;
		    ms <= ms_511;
		end
		ms_511: begin
		    q <= 16'h7e0e;
		    ms <= ms_512;
		end
		ms_512: begin
		    q <= 16'h7e0a;
		    ms <= ms_513;
		end
		ms_513: begin
		    q <= 16'h7e07;
		    ms <= ms_514;
		end
		ms_514: begin
		    q <= 16'h7e04;
		    ms <= ms_515;
		end
		ms_515: begin
		    q <= 16'h7e01;
		    ms <= ms_516;
		end
		ms_516: begin
		    q <= 16'h7dfd;
		    ms <= ms_517;
		end
		ms_517: begin
		    q <= 16'h7dfa;
		    ms <= ms_518;
		end
		ms_518: begin
		    q <= 16'h7df7;
		    ms <= ms_519;
		end
		ms_519: begin
		    q <= 16'h7df4;
		    ms <= ms_520;
		end
		ms_520: begin
		    q <= 16'h7df1;
		    ms <= ms_521;
		end
		ms_521: begin
		    q <= 16'h7dee;
		    ms <= ms_522;
		end
		ms_522: begin
		    q <= 16'h7deb;
		    ms <= ms_523;
		end
		ms_523: begin
		    q <= 16'h7de8;
		    ms <= ms_524;
		end
		ms_524: begin
		    q <= 16'h7de5;
		    ms <= ms_525;
		end
		ms_525: begin
		    q <= 16'h7de2;
		    ms <= ms_526;
		end
		ms_526: begin
		    q <= 16'h7ddf;
		    ms <= ms_527;
		end
		ms_527: begin
		    q <= 16'h7ddc;
		    ms <= ms_528;
		end
		ms_528: begin
		    q <= 16'h7dd9;
		    ms <= ms_529;
		end
		ms_529: begin
		    q <= 16'h7dd7;
		    ms <= ms_530;
		end
		ms_530: begin
		    q <= 16'h7dd4;
		    ms <= ms_531;
		end
		ms_531: begin
		    q <= 16'h7dd1;
		    ms <= ms_532;
		end
		ms_532: begin
		    q <= 16'h7dcf;
		    ms <= ms_533;
		end
		ms_533: begin
		    q <= 16'h7dcc;
		    ms <= ms_534;
		end
		ms_534: begin
		    q <= 16'h7dc9;
		    ms <= ms_535;
		end
		ms_535: begin
		    q <= 16'h7dc7;
		    ms <= ms_536;
		end
		ms_536: begin
		    q <= 16'h7dc4;
		    ms <= ms_537;
		end
		ms_537: begin
		    q <= 16'h7dc2;
		    ms <= ms_538;
		end
		ms_538: begin
		    q <= 16'h7dbf;
		    ms <= ms_539;
		end
		ms_539: begin
		    q <= 16'h7dbd;
		    ms <= ms_540;
		end
		ms_540: begin
		    q <= 16'h7dba;
		    ms <= ms_541;
		end
		ms_541: begin
		    q <= 16'h7db8;
		    ms <= ms_542;
		end
		ms_542: begin
		    q <= 16'h7db6;
		    ms <= ms_543;
		end
		ms_543: begin
		    q <= 16'h7db3;
		    ms <= ms_544;
		end
		ms_544: begin
		    q <= 16'h7db1;
		    ms <= ms_545;
		end
		ms_545: begin
		    q <= 16'h7daf;
		    ms <= ms_546;
		end
		ms_546: begin
		    q <= 16'h7dad;
		    ms <= ms_547;
		end
		ms_547: begin
		    q <= 16'h7dab;
		    ms <= ms_548;
		end
		ms_548: begin
		    q <= 16'h7da9;
		    ms <= ms_549;
		end
		ms_549: begin
		    q <= 16'h7da7;
		    ms <= ms_550;
		end
		ms_550: begin
		    q <= 16'h7da5;
		    ms <= ms_551;
		end
		ms_551: begin
		    q <= 16'h7da3;
		    ms <= ms_552;
		end
		ms_552: begin
		    q <= 16'h7da1;
		    ms <= ms_553;
		end
		ms_553: begin
		    q <= 16'h7d9f;
		    ms <= ms_554;
		end
		ms_554: begin
		    q <= 16'h7d9d;
		    ms <= ms_555;
		end
		ms_555: begin
		    q <= 16'h7d9b;
		    ms <= ms_556;
		end
		ms_556: begin
		    q <= 16'h7d99;
		    ms <= ms_557;
		end
		ms_557: begin
		    q <= 16'h7d97;
		    ms <= ms_558;
		end
		ms_558: begin
		    q <= 16'h7d96;
		    ms <= ms_559;
		end
		ms_559: begin
		    q <= 16'h7d94;
		    ms <= ms_560;
		end
		ms_560: begin
		    q <= 16'h7d92;
		    ms <= ms_561;
		end
		ms_561: begin
		    q <= 16'h7d91;
		    ms <= ms_562;
		end
		ms_562: begin
		    q <= 16'h7d8f;
		    ms <= ms_563;
		end
		ms_563: begin
		    q <= 16'h7d8e;
		    ms <= ms_564;
		end
		ms_564: begin
		    q <= 16'h7d8c;
		    ms <= ms_565;
		end
		ms_565: begin
		    q <= 16'h7d8b;
		    ms <= ms_566;
		end
		ms_566: begin
		    q <= 16'h7d89;
		    ms <= ms_567;
		end
		ms_567: begin
		    q <= 16'h7d88;
		    ms <= ms_568;
		end
		ms_568: begin
		    q <= 16'h7d87;
		    ms <= ms_569;
		end
		ms_569: begin
		    q <= 16'h7d85;
		    ms <= ms_570;
		end
		ms_570: begin
		    q <= 16'h7d84;
		    ms <= ms_571;
		end
		ms_571: begin
		    q <= 16'h7d83;
		    ms <= ms_572;
		end
		ms_572: begin
		    q <= 16'h7d82;
		    ms <= ms_573;
		end
		ms_573: begin
		    q <= 16'h7d80;
		    ms <= ms_574;
		end
		ms_574: begin
		    q <= 16'h7d7f;
		    ms <= ms_575;
		end
		ms_575: begin
		    q <= 16'h7d7e;
		    ms <= ms_576;
		end
		ms_576: begin
		    q <= 16'h7d7d;
		    ms <= ms_577;
		end
		ms_577: begin
		    q <= 16'h7d7c;
		    ms <= ms_578;
		end
		ms_578: begin
		    q <= 16'h7d7b;
		    ms <= ms_579;
		end
		ms_579: begin
		    q <= 16'h7d7a;
		    ms <= ms_580;
		end
		ms_580: begin
		    q <= 16'h7d7a;
		    ms <= ms_581;
		end
		ms_581: begin
		    q <= 16'h7d79;
		    ms <= ms_582;
		end
		ms_582: begin
		    q <= 16'h7d78;
		    ms <= ms_583;
		end
		ms_583: begin
		    q <= 16'h7d77;
		    ms <= ms_584;
		end
		ms_584: begin
		    q <= 16'h7d76;
		    ms <= ms_585;
		end
		ms_585: begin
		    q <= 16'h7d76;
		    ms <= ms_586;
		end
		ms_586: begin
		    q <= 16'h7d75;
		    ms <= ms_587;
		end
		ms_587: begin
		    q <= 16'h7d75;
		    ms <= ms_588;
		end
		ms_588: begin
		    q <= 16'h7d74;
		    ms <= ms_589;
		end
		ms_589: begin
		    q <= 16'h7d74;
		    ms <= ms_590;
		end
		ms_590: begin
		    q <= 16'h7d73;
		    ms <= ms_591;
		end
		ms_591: begin
		    q <= 16'h7d73;
		    ms <= ms_592;
		end
		ms_592: begin
		    q <= 16'h7d72;
		    ms <= ms_593;
		end
		ms_593: begin
		    q <= 16'h7d72;
		    ms <= ms_594;
		end
		ms_594: begin
		    q <= 16'h7d72;
		    ms <= ms_595;
		end
		ms_595: begin
		    q <= 16'h7d71;
		    ms <= ms_596;
		end
		ms_596: begin
		    q <= 16'h7d71;
		    ms <= ms_597;
		end
		ms_597: begin
		    q <= 16'h7d71;
		    ms <= ms_598;
		end
		ms_598: begin
		    q <= 16'h7d71;
		    ms <= ms_599;
		end
		ms_599: begin
		    q <= 16'h7d71;
		    ms <= ms_600;
		end
		ms_600: begin
		    q <= 16'h7d71;
		    ms <= ms_601;
		end
		ms_601: begin
		    q <= 16'h7d71;
		    ms <= ms_602;
		end
		ms_602: begin
		    q <= 16'h7d71;
		    ms <= ms_603;
		end
		ms_603: begin
		    q <= 16'h7d71;
		    ms <= ms_604;
		end
		ms_604: begin
		    q <= 16'h7d71;
		    ms <= ms_605;
		end
		ms_605: begin
		    q <= 16'h7d71;
		    ms <= ms_606;
		end
		ms_606: begin
		    q <= 16'h7d71;
		    ms <= ms_607;
		end
		ms_607: begin
		    q <= 16'h7d71;
		    ms <= ms_608;
		end
		ms_608: begin
		    q <= 16'h7d72;
		    ms <= ms_609;
		end
		ms_609: begin
		    q <= 16'h7d72;
		    ms <= ms_610;
		end
		ms_610: begin
		    q <= 16'h7d72;
		    ms <= ms_611;
		end
		ms_611: begin
		    q <= 16'h7d73;
		    ms <= ms_612;
		end
		ms_612: begin
		    q <= 16'h7d73;
		    ms <= ms_613;
		end
		ms_613: begin
		    q <= 16'h7d74;
		    ms <= ms_614;
		end
		ms_614: begin
		    q <= 16'h7d74;
		    ms <= ms_615;
		end
		ms_615: begin
		    q <= 16'h7d75;
		    ms <= ms_616;
		end
		ms_616: begin
		    q <= 16'h7d75;
		    ms <= ms_617;
		end
		ms_617: begin
		    q <= 16'h7d76;
		    ms <= ms_618;
		end
		ms_618: begin
		    q <= 16'h7d76;
		    ms <= ms_619;
		end
		ms_619: begin
		    q <= 16'h7d77;
		    ms <= ms_620;
		end
		ms_620: begin
		    q <= 16'h7d78;
		    ms <= ms_621;
		end
		ms_621: begin
		    q <= 16'h7d79;
		    ms <= ms_622;
		end
		ms_622: begin
		    q <= 16'h7d7a;
		    ms <= ms_623;
		end
		ms_623: begin
		    q <= 16'h7d7a;
		    ms <= ms_624;
		end
		ms_624: begin
		    q <= 16'h7d7b;
		    ms <= ms_625;
		end
		ms_625: begin
		    q <= 16'h7d7c;
		    ms <= ms_626;
		end
		ms_626: begin
		    q <= 16'h7d7d;
		    ms <= ms_627;
		end
		ms_627: begin
		    q <= 16'h7d7e;
		    ms <= ms_628;
		end
		ms_628: begin
		    q <= 16'h7d7f;
		    ms <= ms_629;
		end
		ms_629: begin
		    q <= 16'h7d80;
		    ms <= ms_630;
		end
		ms_630: begin
		    q <= 16'h7d82;
		    ms <= ms_631;
		end
		ms_631: begin
		    q <= 16'h7d83;
		    ms <= ms_632;
		end
		ms_632: begin
		    q <= 16'h7d84;
		    ms <= ms_633;
		end
		ms_633: begin
		    q <= 16'h7d85;
		    ms <= ms_634;
		end
		ms_634: begin
		    q <= 16'h7d87;
		    ms <= ms_635;
		end
		ms_635: begin
		    q <= 16'h7d88;
		    ms <= ms_636;
		end
		ms_636: begin
		    q <= 16'h7d89;
		    ms <= ms_637;
		end
		ms_637: begin
		    q <= 16'h7d8b;
		    ms <= ms_638;
		end
		ms_638: begin
		    q <= 16'h7d8c;
		    ms <= ms_639;
		end
		ms_639: begin
		    q <= 16'h7d8e;
		    ms <= ms_640;
		end
		ms_640: begin
		    q <= 16'h7d8f;
		    ms <= ms_641;
		end
		ms_641: begin
		    q <= 16'h7d91;
		    ms <= ms_642;
		end
		ms_642: begin
		    q <= 16'h7d92;
		    ms <= ms_643;
		end
		ms_643: begin
		    q <= 16'h7d94;
		    ms <= ms_644;
		end
		ms_644: begin
		    q <= 16'h7d96;
		    ms <= ms_645;
		end
		ms_645: begin
		    q <= 16'h7d97;
		    ms <= ms_646;
		end
		ms_646: begin
		    q <= 16'h7d99;
		    ms <= ms_647;
		end
		ms_647: begin
		    q <= 16'h7d9b;
		    ms <= ms_648;
		end
		ms_648: begin
		    q <= 16'h7d9d;
		    ms <= ms_649;
		end
		ms_649: begin
		    q <= 16'h7d9f;
		    ms <= ms_650;
		end
		ms_650: begin
		    q <= 16'h7da1;
		    ms <= ms_651;
		end
		ms_651: begin
		    q <= 16'h7da3;
		    ms <= ms_652;
		end
		ms_652: begin
		    q <= 16'h7da5;
		    ms <= ms_653;
		end
		ms_653: begin
		    q <= 16'h7da7;
		    ms <= ms_654;
		end
		ms_654: begin
		    q <= 16'h7da9;
		    ms <= ms_655;
		end
		ms_655: begin
		    q <= 16'h7dab;
		    ms <= ms_656;
		end
		ms_656: begin
		    q <= 16'h7dad;
		    ms <= ms_657;
		end
		ms_657: begin
		    q <= 16'h7daf;
		    ms <= ms_658;
		end
		ms_658: begin
		    q <= 16'h7db1;
		    ms <= ms_659;
		end
		ms_659: begin
		    q <= 16'h7db3;
		    ms <= ms_660;
		end
		ms_660: begin
		    q <= 16'h7db6;
		    ms <= ms_661;
		end
		ms_661: begin
		    q <= 16'h7db8;
		    ms <= ms_662;
		end
		ms_662: begin
		    q <= 16'h7dba;
		    ms <= ms_663;
		end
		ms_663: begin
		    q <= 16'h7dbd;
		    ms <= ms_664;
		end
		ms_664: begin
		    q <= 16'h7dbf;
		    ms <= ms_665;
		end
		ms_665: begin
		    q <= 16'h7dc2;
		    ms <= ms_666;
		end
		ms_666: begin
		    q <= 16'h7dc4;
		    ms <= ms_667;
		end
		ms_667: begin
		    q <= 16'h7dc7;
		    ms <= ms_668;
		end
		ms_668: begin
		    q <= 16'h7dc9;
		    ms <= ms_669;
		end
		ms_669: begin
		    q <= 16'h7dcc;
		    ms <= ms_670;
		end
		ms_670: begin
		    q <= 16'h7dcf;
		    ms <= ms_671;
		end
		ms_671: begin
		    q <= 16'h7dd1;
		    ms <= ms_672;
		end
		ms_672: begin
		    q <= 16'h7dd4;
		    ms <= ms_673;
		end
		ms_673: begin
		    q <= 16'h7dd7;
		    ms <= ms_674;
		end
		ms_674: begin
		    q <= 16'h7dd9;
		    ms <= ms_675;
		end
		ms_675: begin
		    q <= 16'h7ddc;
		    ms <= ms_676;
		end
		ms_676: begin
		    q <= 16'h7ddf;
		    ms <= ms_677;
		end
		ms_677: begin
		    q <= 16'h7de2;
		    ms <= ms_678;
		end
		ms_678: begin
		    q <= 16'h7de5;
		    ms <= ms_679;
		end
		ms_679: begin
		    q <= 16'h7de8;
		    ms <= ms_680;
		end
		ms_680: begin
		    q <= 16'h7deb;
		    ms <= ms_681;
		end
		ms_681: begin
		    q <= 16'h7dee;
		    ms <= ms_682;
		end
		ms_682: begin
		    q <= 16'h7df1;
		    ms <= ms_683;
		end
		ms_683: begin
		    q <= 16'h7df4;
		    ms <= ms_684;
		end
		ms_684: begin
		    q <= 16'h7df7;
		    ms <= ms_685;
		end
		ms_685: begin
		    q <= 16'h7dfa;
		    ms <= ms_686;
		end
		ms_686: begin
		    q <= 16'h7dfd;
		    ms <= ms_687;
		end
		ms_687: begin
		    q <= 16'h7e01;
		    ms <= ms_688;
		end
		ms_688: begin
		    q <= 16'h7e04;
		    ms <= ms_689;
		end
		ms_689: begin
		    q <= 16'h7e07;
		    ms <= ms_690;
		end
		ms_690: begin
		    q <= 16'h7e0a;
		    ms <= ms_691;
		end
		ms_691: begin
		    q <= 16'h7e0e;
		    ms <= ms_692;
		end
		ms_692: begin
		    q <= 16'h7e11;
		    ms <= ms_693;
		end
		ms_693: begin
		    q <= 16'h7e14;
		    ms <= ms_694;
		end
		ms_694: begin
		    q <= 16'h7e18;
		    ms <= ms_695;
		end
		ms_695: begin
		    q <= 16'h7e1b;
		    ms <= ms_696;
		end
		ms_696: begin
		    q <= 16'h7e1f;
		    ms <= ms_697;
		end
		ms_697: begin
		    q <= 16'h7e22;
		    ms <= ms_698;
		end
		ms_698: begin
		    q <= 16'h7e26;
		    ms <= ms_699;
		end
		ms_699: begin
		    q <= 16'h7e29;
		    ms <= ms_700;
		end
		ms_700: begin
		    q <= 16'h7e2d;
		    ms <= ms_701;
		end
		ms_701: begin
		    q <= 16'h7e31;
		    ms <= ms_702;
		end
		ms_702: begin
		    q <= 16'h7e34;
		    ms <= ms_703;
		end
		ms_703: begin
		    q <= 16'h7e38;
		    ms <= ms_704;
		end
		ms_704: begin
		    q <= 16'h7e3c;
		    ms <= ms_705;
		end
		ms_705: begin
		    q <= 16'h7e3f;
		    ms <= ms_706;
		end
		ms_706: begin
		    q <= 16'h7e43;
		    ms <= ms_707;
		end
		ms_707: begin
		    q <= 16'h7e47;
		    ms <= ms_708;
		end
		ms_708: begin
		    q <= 16'h7e4b;
		    ms <= ms_709;
		end
		ms_709: begin
		    q <= 16'h7e4f;
		    ms <= ms_710;
		end
		ms_710: begin
		    q <= 16'h7e52;
		    ms <= ms_711;
		end
		ms_711: begin
		    q <= 16'h7e56;
		    ms <= ms_712;
		end
		ms_712: begin
		    q <= 16'h7e5a;
		    ms <= ms_713;
		end
		ms_713: begin
		    q <= 16'h7e5e;
		    ms <= ms_714;
		end
		ms_714: begin
		    q <= 16'h7e62;
		    ms <= ms_715;
		end
		ms_715: begin
		    q <= 16'h7e66;
		    ms <= ms_716;
		end
		ms_716: begin
		    q <= 16'h7e6a;
		    ms <= ms_717;
		end
		ms_717: begin
		    q <= 16'h7e6e;
		    ms <= ms_718;
		end
		ms_718: begin
		    q <= 16'h7e72;
		    ms <= ms_719;
		end
		ms_719: begin
		    q <= 16'h7e77;
		    ms <= ms_720;
		end
		ms_720: begin
		    q <= 16'h7e7b;
		    ms <= ms_721;
		end
		ms_721: begin
		    q <= 16'h7e7f;
		    ms <= ms_722;
		end
		ms_722: begin
		    q <= 16'h7e83;
		    ms <= ms_723;
		end
		ms_723: begin
		    q <= 16'h7e87;
		    ms <= ms_724;
		end
		ms_724: begin
		    q <= 16'h7e8b;
		    ms <= ms_725;
		end
		ms_725: begin
		    q <= 16'h7e90;
		    ms <= ms_726;
		end
		ms_726: begin
		    q <= 16'h7e94;
		    ms <= ms_727;
		end
		ms_727: begin
		    q <= 16'h7e98;
		    ms <= ms_728;
		end
		ms_728: begin
		    q <= 16'h7e9d;
		    ms <= ms_729;
		end
		ms_729: begin
		    q <= 16'h7ea1;
		    ms <= ms_730;
		end
		ms_730: begin
		    q <= 16'h7ea5;
		    ms <= ms_731;
		end
		ms_731: begin
		    q <= 16'h7eaa;
		    ms <= ms_732;
		end
		ms_732: begin
		    q <= 16'h7eae;
		    ms <= ms_733;
		end
		ms_733: begin
		    q <= 16'h7eb2;
		    ms <= ms_734;
		end
		ms_734: begin
		    q <= 16'h7eb7;
		    ms <= ms_735;
		end
		ms_735: begin
		    q <= 16'h7ebb;
		    ms <= ms_736;
		end
		ms_736: begin
		    q <= 16'h7ec0;
		    ms <= ms_737;
		end
		ms_737: begin
		    q <= 16'h7ec4;
		    ms <= ms_738;
		end
		ms_738: begin
		    q <= 16'h7ec9;
		    ms <= ms_739;
		end
		ms_739: begin
		    q <= 16'h7ecd;
		    ms <= ms_740;
		end
		ms_740: begin
		    q <= 16'h7ed2;
		    ms <= ms_741;
		end
		ms_741: begin
		    q <= 16'h7ed6;
		    ms <= ms_742;
		end
		ms_742: begin
		    q <= 16'h7edb;
		    ms <= ms_743;
		end
		ms_743: begin
		    q <= 16'h7ee0;
		    ms <= ms_744;
		end
		ms_744: begin
		    q <= 16'h7ee4;
		    ms <= ms_745;
		end
		ms_745: begin
		    q <= 16'h7ee9;
		    ms <= ms_746;
		end
		ms_746: begin
		    q <= 16'h7eee;
		    ms <= ms_747;
		end
		ms_747: begin
		    q <= 16'h7ef2;
		    ms <= ms_748;
		end
		ms_748: begin
		    q <= 16'h7ef7;
		    ms <= ms_749;
		end
		ms_749: begin
		    q <= 16'h7efc;
		    ms <= ms_750;
		end
		ms_750: begin
		    q <= 16'h7f00;
		    ms <= ms_751;
		end
		ms_751: begin
		    q <= 16'h7f05;
		    ms <= ms_752;
		end
		ms_752: begin
		    q <= 16'h7f0a;
		    ms <= ms_753;
		end
		ms_753: begin
		    q <= 16'h7f0f;
		    ms <= ms_754;
		end
		ms_754: begin
		    q <= 16'h7f14;
		    ms <= ms_755;
		end
		ms_755: begin
		    q <= 16'h7f18;
		    ms <= ms_756;
		end
		ms_756: begin
		    q <= 16'h7f1d;
		    ms <= ms_757;
		end
		ms_757: begin
		    q <= 16'h7f22;
		    ms <= ms_758;
		end
		ms_758: begin
		    q <= 16'h7f27;
		    ms <= ms_759;
		end
		ms_759: begin
		    q <= 16'h7f2c;
		    ms <= ms_760;
		end
		ms_760: begin
		    q <= 16'h7f31;
		    ms <= ms_761;
		end
		ms_761: begin
		    q <= 16'h7f35;
		    ms <= ms_762;
		end
		ms_762: begin
		    q <= 16'h7f3a;
		    ms <= ms_763;
		end
		ms_763: begin
		    q <= 16'h7f3f;
		    ms <= ms_764;
		end
		ms_764: begin
		    q <= 16'h7f44;
		    ms <= ms_765;
		end
		ms_765: begin
		    q <= 16'h7f49;
		    ms <= ms_766;
		end
		ms_766: begin
		    q <= 16'h7f4e;
		    ms <= ms_767;
		end
		ms_767: begin
		    q <= 16'h7f53;
		    ms <= ms_768;
		end
		ms_768: begin
		    q <= 16'h7f58;
		    ms <= ms_769;
		end
		ms_769: begin
		    q <= 16'h7f5d;
		    ms <= ms_770;
		end
		ms_770: begin
		    q <= 16'h7f62;
		    ms <= ms_771;
		end
		ms_771: begin
		    q <= 16'h7f67;
		    ms <= ms_772;
		end
		ms_772: begin
		    q <= 16'h7f6c;
		    ms <= ms_773;
		end
		ms_773: begin
		    q <= 16'h7f71;
		    ms <= ms_774;
		end
		ms_774: begin
		    q <= 16'h7f76;
		    ms <= ms_775;
		end
		ms_775: begin
		    q <= 16'h7f7b;
		    ms <= ms_776;
		end
		ms_776: begin
		    q <= 16'h7f80;
		    ms <= ms_777;
		end
		ms_777: begin
		    q <= 16'h7f85;
		    ms <= ms_778;
		end
		ms_778: begin
		    q <= 16'h7f8a;
		    ms <= ms_779;
		end
		ms_779: begin
		    q <= 16'h7f8f;
		    ms <= ms_780;
		end
		ms_780: begin
		    q <= 16'h7f94;
		    ms <= ms_781;
		end
		ms_781: begin
		    q <= 16'h7f99;
		    ms <= ms_782;
		end
		ms_782: begin
		    q <= 16'h7f9f;
		    ms <= ms_783;
		end
		ms_783: begin
		    q <= 16'h7fa4;
		    ms <= ms_784;
		end
		ms_784: begin
		    q <= 16'h7fa9;
		    ms <= ms_785;
		end
		ms_785: begin
		    q <= 16'h7fae;
		    ms <= ms_786;
		end
		ms_786: begin
		    q <= 16'h7fb3;
		    ms <= ms_787;
		end
		ms_787: begin
		    q <= 16'h7fb8;
		    ms <= ms_788;
		end
		ms_788: begin
		    q <= 16'h7fbd;
		    ms <= ms_789;
		end
		ms_789: begin
		    q <= 16'h7fc2;
		    ms <= ms_790;
		end
		ms_790: begin
		    q <= 16'h7fc7;
		    ms <= ms_791;
		end
		ms_791: begin
		    q <= 16'h7fcd;
		    ms <= ms_792;
		end
		ms_792: begin
		    q <= 16'h7fd2;
		    ms <= ms_793;
		end
		ms_793: begin
		    q <= 16'h7fd7;
		    ms <= ms_794;
		end
		ms_794: begin
		    q <= 16'h7fdc;
		    ms <= ms_795;
		end
		ms_795: begin
		    q <= 16'h7fe1;
		    ms <= ms_796;
		end
		ms_796: begin
		    q <= 16'h7fe6;
		    ms <= ms_797;
		end
		ms_797: begin
		    q <= 16'h7feb;
		    ms <= ms_798;
		end
		ms_798: begin
		    q <= 16'h7ff1;
		    ms <= ms_799;
		end
		ms_799: begin
		    q <= 16'h7ff6;
		    ms <= ms_800;
		end
		ms_800: begin
		    q <= 16'h7ffb;
		    if (send) begin
		        ms <= ms_1;
		    end else begin
		        ms <= ms_pause;
		    end
		end
		default: begin
		    q <= 16'h8000;
		    ms <= ms_pause;
		end
	    endcase
	end
end

endmodule
